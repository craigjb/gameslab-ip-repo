
`timescale 1 ns / 1 ps

	module gslcd_v1_0 #
	(
   		// Parameters of Axi Slave Bus Interface S00_AXI
        parameter integer C_S00_AXI_BASEADDR = 32'h0,
        parameter integer C_S00_AXI_HIGHADDR = 32'h0,
		parameter integer C_S00_AXI_DATA_WIDTH	= 32,
		parameter integer C_S00_AXI_ADDR_WIDTH	= 32,

		// Parameters of Axi Master Bus Interface M00_AXI
		parameter integer C_M00_AXI_BURST_LEN	= 16,
		parameter integer C_M00_AXI_ID_WIDTH	= 1,
		parameter integer C_M00_AXI_ADDR_WIDTH	= 32,
		parameter integer C_M00_AXI_DATA_WIDTH	= 32,
		parameter integer C_M00_AXI_AWUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_ARUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_WUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_RUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_BUSER_WIDTH	= 0
	)
	(
        // Ports of the LCD
        input wire LCD_PCLK,
        output wire LCD_DEN,
        output wire LCD_VSYNC,
        output wire LCD_HSYNC,
        output wire [23 : 0] LCD_DATA,

		// Ports of Axi Slave Bus Interface S00_AXI
        input wire  s00_axi_aclk,
        input wire  s00_axi_aresetn,
        input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
        input wire [2 : 0] s00_axi_awprot,
        input wire  s00_axi_awvalid,
        output wire  s00_axi_awready,
        input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
        input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
        input wire  s00_axi_wvalid,
        output wire  s00_axi_wready,
        output wire [1 : 0] s00_axi_bresp,
        output wire  s00_axi_bvalid,
        input wire  s00_axi_bready,
        input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
        input wire [2 : 0] s00_axi_arprot,
        input wire  s00_axi_arvalid,
        output wire  s00_axi_arready,
        output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
        output wire [1 : 0] s00_axi_rresp,
        output wire  s00_axi_rvalid,
        input wire  s00_axi_rready,

		// Ports of Axi Master Bus Interface M00_AXI
        input wire  m00_axi_aclk,
        input wire  m00_axi_aresetn,
        output wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_awid,
        output wire [C_M00_AXI_ADDR_WIDTH-1 : 0] m00_axi_awaddr,
        output wire [7 : 0] m00_axi_awlen,
        output wire [2 : 0] m00_axi_awsize,
        output wire [1 : 0] m00_axi_awburst,
        output wire  m00_axi_awlock,
        output wire [3 : 0] m00_axi_awcache,
        output wire [2 : 0] m00_axi_awprot,
        output wire [3 : 0] m00_axi_awqos,
        output wire [C_M00_AXI_AWUSER_WIDTH-1 : 0] m00_axi_awuser,
        output wire  m00_axi_awvalid,
        input wire  m00_axi_awready,
        output wire [C_M00_AXI_DATA_WIDTH-1 : 0] m00_axi_wdata,
        output wire [C_M00_AXI_DATA_WIDTH/8-1 : 0] m00_axi_wstrb,
        output wire  m00_axi_wlast,
        output wire [C_M00_AXI_WUSER_WIDTH-1 : 0] m00_axi_wuser,
        output wire  m00_axi_wvalid,
        input wire  m00_axi_wready,
        input wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_bid,
        input wire [1 : 0] m00_axi_bresp,
        input wire [C_M00_AXI_BUSER_WIDTH-1 : 0] m00_axi_buser,
        input wire  m00_axi_bvalid,
        output wire  m00_axi_bready,
        output wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_arid,
        output wire [C_M00_AXI_ADDR_WIDTH-1 : 0] m00_axi_araddr,
        output wire [7 : 0] m00_axi_arlen,
        output wire [2 : 0] m00_axi_arsize,
        output wire [1 : 0] m00_axi_arburst,
        output wire  m00_axi_arlock,
        output wire [3 : 0] m00_axi_arcache,
        output wire [2 : 0] m00_axi_arprot,
        output wire [3 : 0] m00_axi_arqos,
        output wire [C_M00_AXI_ARUSER_WIDTH-1 : 0] m00_axi_aruser,
        output wire  m00_axi_arvalid,
        input wire  m00_axi_arready,
        input wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_rid,
        input wire [C_M00_AXI_DATA_WIDTH-1 : 0] m00_axi_rdata,
        input wire [1 : 0] m00_axi_rresp,
        input wire  m00_axi_rlast,
        input wire [C_M00_AXI_RUSER_WIDTH-1 : 0] m00_axi_ruser,
        input wire  m00_axi_rvalid,
        output wire  m00_axi_rready
	);

    wire reset = ~s00_axi_aresetn;
    wire [C_S00_AXI_ADDR_WIDTH - 1 : 0] slave_awaddr = s00_axi_awaddr - C_S00_AXI_BASEADDR;
    wire [C_S00_AXI_ADDR_WIDTH - 1 : 0] slave_araddr = s00_axi_araddr - C_S00_AXI_BASEADDR;

    GSLCD gslcd_impl(
        .clk(s00_axi_aclk),
        .reset(reset),
        .io_slaveBus_aw_valid(s00_axi_awvalid),
        .io_slaveBus_aw_ready(s00_axi_awready),
        .io_slaveBus_aw_payload_addr(slave_awaddr),
        .io_slaveBus_aw_payload_prot(s00_axi_awprot),
        .io_slaveBus_w_valid(s00_axi_wvalid),
        .io_slaveBus_w_ready(s00_axi_wready),
        .io_slaveBus_w_payload_data(s00_axi_wdata),
        .io_slaveBus_w_payload_strb(s00_axi_wstrb),
        .io_slaveBus_b_valid(s00_axi_bvalid),
        .io_slaveBus_b_ready(s00_axi_bready),
        .io_slaveBus_b_payload_resp(s00_axi_bresp),
        .io_slaveBus_ar_valid(s00_axi_arvalid),
        .io_slaveBus_ar_ready(s00_axi_arready),
        .io_slaveBus_ar_payload_addr(slave_araddr),
        .io_slaveBus_ar_payload_prot(s00_axi_arprot),
        .io_slaveBus_r_valid(s00_axi_rvalid),
        .io_slaveBus_r_ready(s00_axi_rready),
        .io_slaveBus_r_payload_data(s00_axi_rdata),
        .io_slaveBus_r_payload_resp(s00_axi_rresp),
        .io_pclk(LCD_PCLK),
        .io_den(LCD_DEN),
        .io_vsync(LCD_VSYNC),
        .io_hsync(LCD_HSYNC),
        .io_data(LCD_DATA)
    );

	endmodule
