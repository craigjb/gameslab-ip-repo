
`timescale 1 ns / 1 ps

	module gslcd_v1_0 #
	(
        // Parameters for the LCD
        parameter integer C_FRAME_WIDTH = 800,
        parameter integer C_FRAME_HEIGHT = 480,
        parameter integer C_LCD_LINE_REG_WIDTH = 10,
        parameter integer C_LCD_PIXEL_REG_WIDTH = 10,
        parameter integer C_LCD_LINES = 525,
        parameter integer C_LCD_VSYNC_START = 13,
        parameter integer C_LCD_VSYNC_END = 16,
        parameter integer C_LCD_VACTIVE_START = 45,
        parameter integer C_LCD_HPIXELS = 928,
        parameter integer C_LCD_HSYNC_START = 40,
        parameter integer C_LCD_HSYNC_END = 88,
        parameter integer C_LCD_HACTIVE_START = 128,

		// Parameters of Axi Slave Bus Interface S00_AXI
		parameter integer C_S00_AXI_DATA_WIDTH	= 32,
		parameter integer C_S00_AXI_ADDR_WIDTH	= 4,

		// Parameters of Axi Master Bus Interface M00_AXI
		parameter integer C_M00_AXI_BURST_LEN	= 16,
		parameter integer C_M00_AXI_ID_WIDTH	= 1,
		parameter integer C_M00_AXI_ADDR_WIDTH	= 32,
		parameter integer C_M00_AXI_DATA_WIDTH	= 32,
		parameter integer C_M00_AXI_AWUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_ARUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_WUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_RUSER_WIDTH	= 0,
		parameter integer C_M00_AXI_BUSER_WIDTH	= 0
	)
	(
        // Ports of the LCD
        input wire LCD_PCLK,
        output wire LCD_DEN,
        output wire LCD_VSYNC,
        output wire LCD_HSYNC,
        output wire [23 : 0] LCD_DATA,

		// Ports of Axi Slave Bus Interface S00_AXI
        input wire  s00_axi_aclk,
        input wire  s00_axi_aresetn,
        input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
        input wire [2 : 0] s00_axi_awprot,
        input wire  s00_axi_awvalid,
        output wire  s00_axi_awready,
        input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
        input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
        input wire  s00_axi_wvalid,
        output wire  s00_axi_wready,
        output wire [1 : 0] s00_axi_bresp,
        output wire  s00_axi_bvalid,
        input wire  s00_axi_bready,
        input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
        input wire [2 : 0] s00_axi_arprot,
        input wire  s00_axi_arvalid,
        output wire  s00_axi_arready,
        output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
        output wire [1 : 0] s00_axi_rresp,
        output wire  s00_axi_rvalid,
        input wire  s00_axi_rready,

		// Ports of Axi Master Bus Interface M00_AXI
        input wire  m00_axi_aclk,
        input wire  m00_axi_aresetn,
        output wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_awid,
        output wire [C_M00_AXI_ADDR_WIDTH-1 : 0] m00_axi_awaddr,
        output wire [7 : 0] m00_axi_awlen,
        output wire [2 : 0] m00_axi_awsize,
        output wire [1 : 0] m00_axi_awburst,
        output wire  m00_axi_awlock,
        output wire [3 : 0] m00_axi_awcache,
        output wire [2 : 0] m00_axi_awprot,
        output wire [3 : 0] m00_axi_awqos,
        output wire [C_M00_AXI_AWUSER_WIDTH-1 : 0] m00_axi_awuser,
        output wire  m00_axi_awvalid,
        input wire  m00_axi_awready,
        output wire [C_M00_AXI_DATA_WIDTH-1 : 0] m00_axi_wdata,
        output wire [C_M00_AXI_DATA_WIDTH/8-1 : 0] m00_axi_wstrb,
        output wire  m00_axi_wlast,
        output wire [C_M00_AXI_WUSER_WIDTH-1 : 0] m00_axi_wuser,
        output wire  m00_axi_wvalid,
        input wire  m00_axi_wready,
        input wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_bid,
        input wire [1 : 0] m00_axi_bresp,
        input wire [C_M00_AXI_BUSER_WIDTH-1 : 0] m00_axi_buser,
        input wire  m00_axi_bvalid,
        output wire  m00_axi_bready,
        output wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_arid,
        output wire [C_M00_AXI_ADDR_WIDTH-1 : 0] m00_axi_araddr,
        output wire [7 : 0] m00_axi_arlen,
        output wire [2 : 0] m00_axi_arsize,
        output wire [1 : 0] m00_axi_arburst,
        output wire  m00_axi_arlock,
        output wire [3 : 0] m00_axi_arcache,
        output wire [2 : 0] m00_axi_arprot,
        output wire [3 : 0] m00_axi_arqos,
        output wire [C_M00_AXI_ARUSER_WIDTH-1 : 0] m00_axi_aruser,
        output wire  m00_axi_arvalid,
        input wire  m00_axi_arready,
        input wire [C_M00_AXI_ID_WIDTH-1 : 0] m00_axi_rid,
        input wire [C_M00_AXI_DATA_WIDTH-1 : 0] m00_axi_rdata,
        input wire [1 : 0] m00_axi_rresp,
        input wire  m00_axi_rlast,
        input wire [C_M00_AXI_RUSER_WIDTH-1 : 0] m00_axi_ruser,
        input wire  m00_axi_rvalid,
        output wire  m00_axi_rready
	);

    wire lcd_enable;
    wire [C_S00_AXI_DATA_WIDTH-1 : 0] frame_ptr;
    wire active;
    wire rd_active;
    wire frame_start;

    assign LCD_DEN = active;

    gslcd_v1_0_timing # (
      .C_LCD_LINE_REG_WIDTH(C_LCD_LINE_REG_WIDTH),
      .C_LCD_PIXEL_REG_WIDTH(C_LCD_PIXEL_REG_WIDTH),
      .C_LCD_LINES(C_LCD_LINES),
      .C_LCD_VSYNC_START(C_LCD_VSYNC_START),
      .C_LCD_VSYNC_END(C_LCD_VSYNC_END),
      .C_LCD_VACTIVE_START(C_LCD_VACTIVE_START),
      .C_LCD_HPIXELS(C_LCD_HPIXELS),
      .C_LCD_HSYNC_START(C_LCD_HSYNC_START),
      .C_LCD_HSYNC_END(C_LCD_HSYNC_END),
      .C_LCD_HACTIVE_START(C_LCD_HACTIVE_START)
    ) gslcd_v1_0_timing_inst (
      .PCLK(LCD_PCLK),
      .EN(lcd_enable),
      .VSYNC(LCD_VSYNC),
      .HSYNC(LCD_HSYNC),
      .ACTIVE(active),
      .RD_ACTIVE(rd_active),
      .FRAME_START(frame_start)
    );

    // Instantiation of Axi Bus Interface S00_AXI
    gslcd_v1_0_S00_AXI # ( 
        .C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
        .C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH)
    ) gslcd_v1_0_S00_AXI_inst (
        .S_AXI_ACLK(s00_axi_aclk),
        .S_AXI_ARESETN(s00_axi_aresetn),
        .S_AXI_AWADDR(s00_axi_awaddr),
        .S_AXI_AWPROT(s00_axi_awprot),
        .S_AXI_AWVALID(s00_axi_awvalid),
        .S_AXI_AWREADY(s00_axi_awready),
        .S_AXI_WDATA(s00_axi_wdata),
        .S_AXI_WSTRB(s00_axi_wstrb),
        .S_AXI_WVALID(s00_axi_wvalid),
        .S_AXI_WREADY(s00_axi_wready),
        .S_AXI_BRESP(s00_axi_bresp),
        .S_AXI_BVALID(s00_axi_bvalid),
        .S_AXI_BREADY(s00_axi_bready),
        .S_AXI_ARADDR(s00_axi_araddr),
        .S_AXI_ARPROT(s00_axi_arprot),
        .S_AXI_ARVALID(s00_axi_arvalid),
        .S_AXI_ARREADY(s00_axi_arready),
        .S_AXI_RDATA(s00_axi_rdata),
        .S_AXI_RRESP(s00_axi_rresp),
        .S_AXI_RVALID(s00_axi_rvalid),
        .S_AXI_RREADY(s00_axi_rready),
        .LCD_ENABLE(lcd_enable),
        .FRAME_PTR(frame_ptr)
    );

    wire fifo_rst;
    wire [ C_M00_AXI_DATA_WIDTH-1 : 0 ] fifo_din;
    wire fifo_wren;
    wire fifo_almost_full;
    wire fifo_full;
    wire fifo_rden;
    wire fifo_empty;
    wire [ C_M00_AXI_DATA_WIDTH-1 : 0 ] fifo_dout;

    FIFO36 # (
        .DATA_WIDTH(36),
        .ALMOST_FULL_OFFSET(13'h10),
        .ALMOST_EMPTY_OFFSET(13'h10)
    ) fifo_inst (
        .DI(fifo_din),
        .WREN(fifo_wren),
        .WRCLK(m00_axi_aclk),
        .RST(fifo_rst),
        .ALMOSTFULL(fifo_almost_full),
        .FULL(fifo_full),
        .RDCLK(LCD_PCLK),
        .RDEN(fifo_rden),
        .DO(fifo_dout),
        .EMPTY(fifo_empty)
    );

    wire [ 23 : 0 ]data24;

    gslcd_v1_0_fifo_32to24 fifo_32to24_inst (
        .clk(LCD_PCLK),
        .reset(FRAME_START),
        .rd_en(rd_active),
        .data32(fifo_dout),
        .data24(data24),
        .rd_en32(fifo_rden)
    );

    assign LCD_DATA = fifo_empty ? 24'hff0000 : data24;

    //// Instantiation of Axi Bus Interface M00_AXI
    gslcd_v1_0_M00_AXI # ( 
        .C_M_AXI_BURST_LEN(C_M00_AXI_BURST_LEN),
        .C_M_AXI_ID_WIDTH(C_M00_AXI_ID_WIDTH),
        .C_M_AXI_ADDR_WIDTH(C_M00_AXI_ADDR_WIDTH),
        .C_M_AXI_DATA_WIDTH(C_M00_AXI_DATA_WIDTH),
        .C_M_AXI_AWUSER_WIDTH(C_M00_AXI_AWUSER_WIDTH),
        .C_M_AXI_ARUSER_WIDTH(C_M00_AXI_ARUSER_WIDTH),
        .C_M_AXI_WUSER_WIDTH(C_M00_AXI_WUSER_WIDTH),
        .C_M_AXI_RUSER_WIDTH(C_M00_AXI_RUSER_WIDTH),
        .C_M_AXI_BUSER_WIDTH(C_M00_AXI_BUSER_WIDTH),
        .C_LCD_DATA_LEN(C_FRAME_WIDTH * C_FRAME_HEIGHT * 3)
    ) gslcd_v1_0_M00_AXI_inst (
        .M_AXI_ACLK(m00_axi_aclk),
        .M_AXI_ARESETN(m00_axi_aresetn),
        .M_AXI_AWID(m00_axi_awid),
        .M_AXI_AWADDR(m00_axi_awaddr),
        .M_AXI_AWLEN(m00_axi_awlen),
        .M_AXI_AWSIZE(m00_axi_awsize),
        .M_AXI_AWBURST(m00_axi_awburst),
        .M_AXI_AWLOCK(m00_axi_awlock),
        .M_AXI_AWCACHE(m00_axi_awcache),
        .M_AXI_AWPROT(m00_axi_awprot),
        .M_AXI_AWQOS(m00_axi_awqos),
        .M_AXI_AWUSER(m00_axi_awuser),
        .M_AXI_AWVALID(m00_axi_awvalid),
        .M_AXI_AWREADY(m00_axi_awready),
        .M_AXI_WDATA(m00_axi_wdata),
        .M_AXI_WSTRB(m00_axi_wstrb),
        .M_AXI_WLAST(m00_axi_wlast),
        .M_AXI_WUSER(m00_axi_wuser),
        .M_AXI_WVALID(m00_axi_wvalid),
        .M_AXI_WREADY(m00_axi_wready),
        .M_AXI_BID(m00_axi_bid),
        .M_AXI_BRESP(m00_axi_bresp),
        .M_AXI_BUSER(m00_axi_buser),
        .M_AXI_BVALID(m00_axi_bvalid),
        .M_AXI_BREADY(m00_axi_bready),
        .M_AXI_ARID(m00_axi_arid),
        .M_AXI_ARADDR(m00_axi_araddr),
        .M_AXI_ARLEN(m00_axi_arlen),
        .M_AXI_ARSIZE(m00_axi_arsize),
        .M_AXI_ARBURST(m00_axi_arburst),
        .M_AXI_ARLOCK(m00_axi_arlock),
        .M_AXI_ARCACHE(m00_axi_arcache),
        .M_AXI_ARPROT(m00_axi_arprot),
        .M_AXI_ARQOS(m00_axi_arqos),
        .M_AXI_ARUSER(m00_axi_aruser),
        .M_AXI_ARVALID(m00_axi_arvalid),
        .M_AXI_ARREADY(m00_axi_arready),
        .M_AXI_RID(m00_axi_rid),
        .M_AXI_RDATA(m00_axi_rdata),
        .M_AXI_RRESP(m00_axi_rresp),
        .M_AXI_RLAST(m00_axi_rlast),
        .M_AXI_RUSER(m00_axi_ruser),
        .M_AXI_RVALID(m00_axi_rvalid),
        .M_AXI_RREADY(m00_axi_rready),
        .FRAME_PTR(frame_ptr),
        .FRAME_START(frame_start),
        .FIFO_RST(fifo_rst),
        .FIFO_DIN(fifo_din),
        .FIFO_WREN(fifo_wren),
        .FIFO_ALMOST_FULL(fifo_almost_full),
        .FIFO_FULL(fifo_full)
    );

	endmodule
